module vcordium

import lib

pub const (
	version = '0.0.0'
)